
module master_controller();




endmodule